 module vraylib


const (
	albedo			= 0
	diffuse			= 0
	metalness		= 1
	normal			= 2
	roughness		= 4
	occlusion		= 5
	emission 		= 6
	height			= 7
	cubemap			= 8
	irradiance		= 9
	prefilter		= 10
	brdf			= 11
)
