module vraylib

// TODO: put here maybe comments/instructions