module vraylib

// --------------------------------------------------------
//  Module: Shapes
// --------------------------------------------------------

fn C.DrawPixel(posX, posY int, color C.Color)
fn C.DrawPixelV(position C.Vector2, color C.Color)
fn C.DrawLine(startPosX, startPosY, endPosX, endPosY int, color C.Color)
fn C.DrawLineV(startPos, endPos C.Vector2, color C.Color)
fn C.DrawLineEx(startPos, endPos C.Vector2, thick f32, color C.Color)
fn C.DrawLineBezier(startPos, endPos C.Vector2, thick f32, color C.Color)
fn C.DrawLineStrip(points C.Vector2, numPoints int, color C.Color)
fn C.DrawCircle(centerX, centerY int, radius f32, color C.Color)
fn C.DrawCircleSector(center C.Vector2, radius f32, startAngle, endAngle, segments int, color C.Color)
fn C.DrawCircleSectorLines(center C.Vector2, radius f32, startAngle, endAngle, segments int, color C.Color)
fn C.DrawCircleGradient(centerX, centerY int, radius f32, coor1, color2 C.Color)
fn C.DrawCircleV(center C.Vector2, radius f32, color C.Color)
fn C.DrawCircleLines(centerX, centerY int, radius f32, color C.Color)
fn C.DrawRing(center C.Vector2, innerRadius, outerRadius f32, startAngle, endAngle, segments int, color C.Color)
fn C.DrawRingLines(center C.Vector2, innerRadius, outerRadius f32, startAngle, endAngle, segments int, color C.Color)
fn C.DrawRectangle(posX, posY, width, height int, color C.Color)
fn C.DrawRectangleV(position, size C.Vector2, color C.Color)
fn C.DrawRectangleRec(rec C.Rectangle, color C.Color)
fn C.DrawRectanglePro(rec C.Rectangle, origin C.Vector2, rotation f32, color C.Color)
fn C.DrawRectangleGradientV(posX, posY, width, height int, color1, color2 C.Color)
fn C.DrawRectangleGradientH(posX, posY, width, height int, color1, color2 C.Color)
fn C.DrawRectangleGradientEx(rec C.Rectangle, col1, col2, col3, col4 C.Color)
fn C.DrawRectangleLines(posX, posY, width, height int, color C.Color)
fn C.DrawRectangleLinesEx(rec C.Rectangle, lineThick int, color C.Color)
fn C.DrawRectangleRounded(rec C.Rectangle, roundness f32, segments int, color C.Color)
fn C.DrawRectangleRoundedLines(rec C.Rectangle, roundness f32, segments, lineThick int, color C.Color)
fn C.DrawTriangle(v1, v2, v3 C.Vector2, color C.Color)
fn C.DrawTriangleLines(v1, v2, v3 C.Vector2, color C.Color)
fn C.DrawTriangleFan(points C.Vector2, numPoints int, color C.Color)
fn C.DrawPoly(center C.Vector2, sides int, radius, rotation f32, color C.Color)

fn C.SetShapesTexture(texture C.Texture2D, source C.Rectangle)

fn C.CheckCollisionRecs(rec1, rec2 C.Rectangle) bool
fn C.CheckCollisionCircles(center1 C.Vector2, radius1 f32, center2 C.Vector2, radius2 f32) bool
fn C.CheckCollisionCircleRec(center C.Vector2, radius f32, rec C.Rectangle) bool
fn C.GetCollisionRec(rec1, rec2 C.Rectangle) C.Rectangle
fn C.CheckCollisionPointRec(point C.Vector2, rec C.Rectangle) bool
fn C.CheckCollisionPointCircle(point C.Vector2, center C.Vector2, radius f32) bool
fn C.CheckCollisionPointTriangle(point, p1, p2, p3 C.Vector3) bool

// Shape Drawing Functions
// Basic shapes drawing functions
pub fn draw_pixel(posX, posY int, color Color) {
	C.DrawPixel(posX, posY, color)
}

pub fn draw_pixel_v(position Vector2, color Color) {
	C.DrawPixelV(position, color)
}

pub fn draw_line(startPosX, startPosY, endPosX, endPosY int, color Color) {
	C.DrawLine(startPosX, startPosY, endPosX, endPosY, color)
}

pub fn draw_line_v(startPos, endPos Vector2, color Color) {
	C.DrawLineV(startPos, endPos, color)
}

pub fn draw_line_ex(startPos, endPos Vector2, thick f32, color Color) {
	C.DrawLineEx(startPos, endPos, thick, color)
}

pub fn draw_line_bezier(startPos, endPos Vector2, thick f32, color Color) {
	C.DrawLineBezier(startPos, endPos, thick, color)
}

pub fn draw_line_strip(points &Vector2, numPoints int, color Color) {
	C.DrawLineStrip(points, numPoints, color)
}

pub fn draw_circle(centerX, centerY int, radius f32, color Color) {
	C.DrawCircle(centerX, centerY, radius, color)
}

pub fn draw_circle_sector(center Vector2, radius f32, startAngle, endAngle, segments int, color Color) {
	C.DrawCircleSector(center, radius, startAngle, endAngle, segments, color)
}

pub fn draw_circle_sector_lines(center Vector2, radius f32, startAngle, endAngle, segments int, color Color) {
	C.DrawCircleSectorLines(center, radius, startAngle, endAngle, segments, color)
}

pub fn draw_circle_gradient(centerX, centerY int, radius f32, color1, color2 Color) {
	C.DrawCircleGradient(centerX, centerY, radius, color1, color2)
}

pub fn draw_circle_v(center Vector2, radius f32, color Color) {
	C.DrawCircleV(center, radius, color)
}

pub fn draw_circle_lines(centerX, centerY int, radius f32, color Color) {
	C.DrawCircleLines(centerX, centerY, radius, color)
}

pub fn draw_ring(center Vector2, innerRadius, outerRadius f32, startAngle, endAngle, segments int, color Color) {
	C.DrawRing(center, innerRadius, outerRadius, startAngle, endAngle, segments, color)
}

pub fn draw_ring_lines(center Vector2, innerRadius, outerRadius f32, startAngle, endAngle, segments int, color Color) {
	C.DrawRingLines(center, innerRadius, outerRadius, startAngle, endAngle, segments, color)
}

pub fn draw_rectangle(posX, posY, width, height int, color Color) {
	C.DrawRectangle(posX, posY, width, height, color)
}

pub fn draw_rectangle_v(position, size Vector2, color Color) {
	C.DrawRectangleV(position, size, color)
}

pub fn draw_rectangle_rec(rec Rectangle, color Color) {
	C.DrawRectangleRec(rec, color)
}

pub fn draw_rectangle_pro(rec Rectangle, origin Vector2, rotation f32, color Color) {
	C.DrawRectanglePro(rec, origin, rotation, color)
}

pub fn draw_rectangle_gradient_v(posX, posY, width, height int, color1, color2 Color) {
	C.DrawRectangleGradientV(posX, posY, width, height, color1, color2)
}

pub fn draw_rectangle_gradient_h(posX, posY, width, height int, color1, color2 Color) {
	C.DrawRectangleGradientH(posX, posY, width, height, color1, color2)
}

pub fn draw_rectangle_gradient_ex(rec Rectangle, col1, col2, col3, col4 Color) {
	C.DrawRectangleGradientEx(rec, col1, col2, col3, col4)
}

pub fn draw_rectangle_lines(posX, posY, width, height int, color Color) {
	C.DrawRectangleLines(posX, posY, width, height, color)
}

pub fn draw_rectangle_lines_ex(rec Rectangle, lineThick int, color Color) {
	C.DrawRectangleLinesEx(rec, lineThick, color)
}

pub fn draw_rectangle_rounded(rec Rectangle, roundness f32, segments int, color Color) {
	C.DrawRectangleRounded(rec, roundness, segments, color)
}

pub fn draw_rectangle_rounded_lines(rec Rectangle, roundness f32, segments, lineThick int, color Color) {
	C.DrawRectangleRoundedLines(rec, roundness, segments, lineThick, color)
}

pub fn draw_triangle(v1, v2, v3 Vector2, color Color) {
	C.DrawTriangle(v1, v2, v3, color)
}

pub fn draw_triangle_lines(v1, v2, v3 Vector2, color Color) {
	C.DrawTriangleLines(v1, v2, v3, color)
}

pub fn draw_triangle_fan(points &Vector2, numPoints int, color Color) {
	C.DrawTriangleFan(points, numPoints, color)
}

pub fn draw_poly(center Vector2, sides int, radius, rotation f32, color Color) {
	C.DrawPoly(center, sides, radius, rotation, color)
}

pub fn set_shapes_texture(texture Texture2D, source Rectangle) {
	C.SetShapesTexture(texture, source)
}

// Basic Shapes Collision Detection Functions
pub fn check_collision_recs(rec1, rec2 Rectangle) bool {
	return C.CheckCollisionRecs(rec1, rec2)
}

pub fn check_collision_circles(center1 Vector2, radius1 f32, center2 Vector2, radius2 f32) bool {
	return C.CheckCollisionCircles(center1, radius1, center2, radius2)
}

pub fn check_collision_circle_rec(center Vector2, radius f32, rec Rectangle) bool {
	return C.CheckCollisionCircleRec(center, radius, rec)
}


pub fn get_collision_rec(rec1, rec2 Rectangle) Rectangle {
	return C.GetCollisionRec(rec1, rec2)
}

pub fn check_collision_point_rec(point Vector2, rec Rectangle) bool {
	return C.CheckCollisionPointRec(point, rec)
}

pub fn check_collision_point_circle(point, center Vector2, radius f32) bool {
	return C.CheckCollisionPointCircle(point, center, radius)
}

pub fn check_collision_point_triangle(point, p1, p2, p3 Vector2) bool {
	return C.CheckCollisionPointTriangle(point, p1, p2, p3)
}

